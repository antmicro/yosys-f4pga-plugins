// Copyright (C) 2022  The SymbiFlow Authors.
//
// Use of this source code is governed by a ISC-style
// license that can be found in the LICENSE file or at
// https://opensource.org/licenses/ISC
//
// SPDX-License-Identifier:ISC

`include "qlf_k6n10f/cells_sim.v"
`timescale 1ns/1ps

`define UPAE1 10
`define UPAF1 10
`define UPAE2 10
`define UPAF2 10
`define SPLIT 0
`define SYNC_FIFO1 0
`define SYNC_FIFO2 0
`define FMODE1 1
`define POWERDN1 0
`define SLEEP1 0
`define PROTECT1 0
`define FMODE2 0
`define POWERDN2 0
`define SLEEP2 0
`define PROTECT2 0
`define RMODE_A1 MODE_36
`define RMODE_B1 MODE_36
`define WMODE_A1 MODE_36
`define WMODE_B1 MODE_36
`define RMODE_A2 MODE_36
`define RMODE_B2 MODE_36
`define WMODE_A2 MODE_36
`define WMODE_B2 MODE_36


module tb;
	localparam W_PERIOD = 30;
	localparam R_PERIOD = 29;
	reg WEN_A1;
	reg WEN_B1;
	reg REN_A1;
	reg REN_B1;
	reg CLK_A1;
	reg CLK_B1;
	reg [1:0] BE_A1;
	reg [1:0] BE_B1;
	reg [14:0] ADDR_A1;
	reg [14:0] ADDR_B1;
	reg [17:0] WDATA_A1;
	reg [17:0] WDATA_B1;
	wire [17:0] RDATA_A1;
	wire [17:0] RDATA_B1;
	wire UNDERRUN1;
	wire OVERRUN1;
	wire UNDERRUN2;
	wire OVERRUN2;
	wire EMPTY1;
	wire EPO1;
	wire EWM1;
	wire FULL1;
	wire FMO1;
	wire FWM1;
	reg FLUSH1;
	reg WEN_A2;
	reg WEN_B2;
	reg REN_A2;
	reg REN_B2;
	reg CLK_A2;
	reg CLK_B2;
	reg [1:0] BE_A2;
	reg [1:0] BE_B2;
	wire [13:0] ADDR_A2;
	wire [13:0] ADDR_B2;
	reg [17:0] WDATA_A2;
	reg [17:0] WDATA_B2;
	wire [17:0] RDATA_A2;
	wire [17:0] RDATA_B2;
	wire EMPTY2;
	wire EPO2;
	wire EWM2;
	wire FULL2;
	wire FMO2;
	wire FWM2;
	reg FLUSH2;
	reg [15:0] RAM_ID_i;
	wire [17:0] RDATA_A18;
	wire [17:0] RDATA_B18;
	wire [8:0] RDATA_A9;
	wire [8:0] RDATA_B9;
	reg PL_INIT_i;
	reg PL_ENA_i;
	reg PL_REN_i;
	reg PL_CLK_i;
	reg [1:0] PL_WEN_i;
	wire [1:0] PL_WEN_o;
	reg [23:0] PL_ADDR_i;
	reg [35:0] PL_DATA_i;
	wire [35:0] PL_DATA_o;
	wire [35:0] expected_data_a;
	wire [35:0] expected_data_b;
	wire [35:0] last_expected_a;
	wire [35:0] last_expected_b;
	wire [17:0] last_expected_a18;
	wire [17:0] last_expected_b18;
	wire [8:0] last_expected_a9;
	wire [8:0] last_expected_b9;
	wire [14:0] last_addr_a;
	wire [14:0] last_addr_b;
	wire valid_a;
	wire valid_b;
	wire [3:0] index4_a;
	wire [3:0] index4_b;
	wire [1:0] index2_a;
	wire [1:0] index2_b;
	wire index_a;
	wire index_b;
	reg last_empty1;
	wire last_empty2;
	wire [35:0] fifo_dout;
	wire [35:0] fifo_din;
	localparam MODE_36 = 3'b011;
	task fA_36x36;
		begin
			$display("%d: Fifo 36-bit write 36-bit read", $time);
			FLUSH1 = 1;
			@(posedge CLK_A1);
			@(posedge CLK_B1);
			FLUSH1 = 0;
		end
	endtask
	task fA_push36;
		input [35:0] data;
		begin
			@(negedge CLK_A1) begin
				WDATA_A2 = data[35:18];
				WDATA_A1 = data[17:0];
				WEN_A1 = 1;
			end
			@(posedge CLK_A1)
				#(2) WEN_A1 = 0;
		end
	endtask
	task fA_pop;
		input [35:0] expected;
		input [35:0] msk;
		begin
			if (last_empty1 || EMPTY1)
				while (EMPTY1 == 1) begin
					@(posedge CLK_B1);
				end
			if (({RDATA_B2, RDATA_B1} & msk) !== expected) begin
				$display("%d: POP FIFO ERROR: mismatch: expected = %9x mask = %5x, actuall = %9x", $time, expected, msk, {RDATA_B2, RDATA_B1});
				error_cnt = error_cnt + 1'b1;
			end
			@(negedge CLK_B1) REN_B1 = 1;
			@(posedge CLK_B1)
				#(2) REN_B1 = 0;
		end
	endtask
	integer wcount_a;
	integer rcount_a;
	integer state_a;
	integer wcount_b;
	integer rcount_b;
	integer state_b;
	integer error_cnt = 0;
	initial CLK_A1 = 0;
	initial CLK_B1 = 0;
	initial CLK_A2 = 0;
	initial CLK_B2 = 0;
	initial forever #(R_PERIOD) CLK_A1 = ~CLK_A1;
	initial forever #(W_PERIOD) CLK_B1 = ~CLK_B1;
	initial forever #(R_PERIOD) CLK_A2 = ~CLK_A2;
	initial forever #(W_PERIOD) CLK_B2 = ~CLK_B2;
	initial begin
		$dumpfile(`VCD_FILE);
		$dumpvars(0, tb);
	end
	initial #(1) begin
		WEN_A1 = 0;
		REN_A1 = 0;
		WEN_B1 = 0;
		REN_B1 = 0;
		BE_A1 = 2'b11;
		BE_A2 = 2'b11;
		BE_B1 = 2'b11;
		BE_B2 = 2'b11;
		ADDR_A1 = 14'b00000000000000;
		ADDR_B1 = 14'b00000000000000;
		WDATA_A1 = 18'b000000000000000000;
		WDATA_B1 = 18'h00000;
		wcount_a = 0;
		rcount_a = 0;
		state_a = 0;
		wcount_b = 0;
		rcount_b = 0;
		state_b = 0;
		PL_INIT_i = 0;
		PL_ADDR_i = 0;
		PL_ENA_i = 0;
		PL_REN_i = 0;
		PL_WEN_i = 2'b00;
		PL_CLK_i = 0;
		PL_DATA_i = 0;
		RAM_ID_i = 16'b0000000000000000;
		WEN_A2 = 0;
		REN_A2 = 0;
		WEN_B2 = 0;
		REN_B2 = 0;
		FLUSH1 = 0;
		FLUSH2 = 0;
	end
	initial begin
		#(100)
		@(posedge CLK_A1);
		@(posedge CLK_B1);
	end
	assign fifo_dout = {RDATA_B2, RDATA_B1};
	assign fifo_din = {WDATA_A2, WDATA_A1};
	assign {EMPTY1, EPO1, EWM1, UNDERRUN1, FULL1, FMO1, FWM1, OVERRUN1} = RDATA_A1[7:0];
	assign {EMPTY2, EPO2, EWM2, UNDERRUN2, FULL2, FMO2, FWM2, OVERRUN2} = RDATA_A2[7:0];
	always @(posedge CLK_B1) last_empty1 <= EMPTY1;
	always @(*)
		case (state_a)
			0: begin
				fA_36x36;
				if (!EMPTY1) begin
					$display("%d: FIFO ERROR: EMPTY flag not set", $time);
					error_cnt = error_cnt + 1'b1;
				end
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				if (!EMPTY1) begin
					$display("%d: FIFO ERROR: EMPTY flag not set", $time);
					error_cnt = error_cnt + 1'b1;
				end
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				if (!EMPTY1) begin
					$display("%d: FIFO ERROR: EMPTY flag not set", $time);
					error_cnt = error_cnt + 1'b1;
				end
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				if (!FULL1) begin
					$display("%d: FIFO ERROR: FULL flag not set", $time);
					error_cnt = error_cnt + 1'b1;
				end
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				if (!EMPTY1) begin
					$display("%d: FIFO ERROR: EMPTY flag not set", $time);
					error_cnt = error_cnt + 1'b1;
				end
				@(posedge CLK_A1);
				@(posedge CLK_B1);
				@(posedge CLK_A1);
				@(posedge CLK_B1);
				@(posedge CLK_A1);
				@(posedge CLK_B1);
				@(posedge CLK_A1);
				@(posedge CLK_B1);
				@(posedge CLK_A1);
				@(posedge CLK_B1);
				@(posedge CLK_A1);
				@(posedge CLK_B1);
				$finish_and_return( (error_cnt == 0) ? 0 : -1 );
			end
		endcase
	wire PL_INIT_o;
	wire PL_ENA_o;
	wire PL_REN_o;
	wire PL_CLK_o;

	TDP36K #(
		.UPAE1_i(`UPAE1),
		.UPAF1_i(`UPAF1),
		.UPAE2_i(`UPAE2),
		.UPAF2_i(`UPAF2),
		.SPLIT_i(`SPLIT),
		.SYNC_FIFO1_i(`SYNC_FIFO1),
		.SYNC_FIFO2_i(`SYNC_FIFO2),
		.FMODE1_i(`FMODE1),
		.POWERDN1_i(`POWERDN1),
		.SLEEP1_i(`SLEEP1),
		.PROTECT1_i(`PROTECT1),
		.FMODE2_i(`FMODE2),
		.POWERDN2_i(`POWERDN2),
		.SLEEP2_i(`SLEEP2),
		.PROTECT2_i(`PROTECT2),
		.RMODE_A1_i(`RMODE_A1),
		.RMODE_B1_i(`RMODE_B1),
		.WMODE_A1_i(`WMODE_A1),
		.WMODE_B1_i(`WMODE_B1),
		.RMODE_A2_i(`RMODE_A2),
		.RMODE_B2_i(`RMODE_B2),
		.WMODE_A2_i(`WMODE_A2),
		.WMODE_B2_i(`WMODE_B2)
	)tdp36_1(
		.CLK_A1_i(CLK_A1),
		.CLK_B1_i(CLK_B1),
		.WEN_A1_i(WEN_A1),
		.WEN_B1_i(WEN_B1),
		.REN_A1_i(REN_A1),
		.REN_B1_i(REN_B1),
		.BE_A1_i(BE_A1),
		.BE_B1_i(BE_B1),
		.ADDR_A1_i(ADDR_A1),
		.ADDR_B1_i(ADDR_B1),
		.WDATA_A1_i(WDATA_A1),
		.WDATA_B1_i(WDATA_B1),
		.RDATA_A1_o(RDATA_A1),
		.RDATA_B1_o(RDATA_B1),
		.FLUSH1_i(FLUSH1),
		.CLK_A2_i(CLK_A2),
		.CLK_B2_i(CLK_B2),
		.WEN_A2_i(WEN_A2),
		.WEN_B2_i(WEN_B2),
		.REN_A2_i(REN_A2),
		.REN_B2_i(REN_B2),
		.BE_A2_i(BE_A2),
		.BE_B2_i(BE_B2),
		.ADDR_A2_i(ADDR_A2),
		.ADDR_B2_i(ADDR_B2),
		.WDATA_A2_i(WDATA_A2),
		.WDATA_B2_i(WDATA_B2),
		.RDATA_A2_o(RDATA_A2),
		.RDATA_B2_o(RDATA_B2),
		.FLUSH2_i(FLUSH2),
		.RAM_ID_i(RAM_ID_i),
		.PL_INIT_i(PL_INIT_i),
		.PL_ENA_i(PL_ENA_i),
		.PL_WEN_i(PL_WEN_i),
		.PL_REN_i(PL_REN_i),
		.PL_CLK_i(PL_CLK_i),
		.PL_ADDR_i(PL_ADDR_i),
		.PL_DATA_i(PL_DATA_i),
		.PL_INIT_o(PL_INIT_o),
		.PL_ENA_o(PL_ENA_o),
		.PL_WEN_o(PL_WEN_o),
		.PL_REN_o(PL_REN_o),
		.PL_CLK_o(PL_CLK_o),
		.PL_ADDR_o(),
		.PL_DATA_o(PL_DATA_o)
	);
endmodule
